`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/03/21 19:08:44
// Design Name: 
// Module Name: MULTU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include "defines.vh"

module MULTU(
    input reset,
    input [`RegBus] a,
    input [`RegBus] b,
    output [`DRegBus] z
    );
    
    reg [`DRegBus] tmp0;
    reg [`DRegBus] tmp1;
    reg [`DRegBus] tmp2;
    reg [`DRegBus] tmp3;
    reg [`DRegBus] tmp4;
    reg [`DRegBus] tmp5;
    reg [`DRegBus] tmp6;
    reg [`DRegBus] tmp7;
    reg [`DRegBus] tmp8;
    reg [`DRegBus] tmp9;
    reg [`DRegBus] tmp10;
    reg [`DRegBus] tmp11;
    reg [`DRegBus] tmp12;
    reg [`DRegBus] tmp13;
    reg [`DRegBus] tmp14;
    reg [`DRegBus] tmp15;
    reg [`DRegBus] tmp16;
    reg [`DRegBus] tmp17;
    reg [`DRegBus] tmp18;
    reg [`DRegBus] tmp19;
    reg [`DRegBus] tmp20;
    reg [`DRegBus] tmp21;
    reg [`DRegBus] tmp22;
    reg [`DRegBus] tmp23;
    reg [`DRegBus] tmp24;
    reg [`DRegBus] tmp25;
    reg [`DRegBus] tmp26;
    reg [`DRegBus] tmp27;
    reg [`DRegBus] tmp28;
    reg [`DRegBus] tmp29;
    reg [`DRegBus] tmp30;
    reg [`DRegBus] tmp31;
    
    wire [`DRegBus] tans_0_1, tans_2_3, tans_4_5, tans_6_7, tans_8_9, tans_10_11, tans_12_13, tans_14_15;
    wire [`DRegBus] tans_16_17, tans_18_19, tans_20_21, tans_22_23, tans_24_25, tans_26_27, tans_28_29, tans_30_31;
    wire [`DRegBus] tans_01_23, tans_45_67, tans_89_1011, tans_1213_1415, tans_1617_1819, tans_2021_2223, tans_2425_2627, tans_2829_3031;
    wire [`DRegBus] tans_0123_4567, tans_891011_12131415, tans_16171819_20212223, tans_24252627_28293031;
    wire [`DRegBus] tans_012345678_9101112131415, tans_1617181920212223_2425262728293031;
    
    assign tans_0_1 = tmp0 + tmp1;
    assign tans_2_3 = tmp2 + tmp3;
    assign tans_4_5 = tmp4 + tmp5;
    assign tans_6_7 = tmp6 + tmp7;
    assign tans_8_9 = tmp8 + tmp9;
    assign tans_10_11 = tmp10 + tmp11;
    assign tans_12_13 = tmp12 + tmp13;
    assign tans_14_15 = tmp14 + tmp15;
    assign tans_16_17 = tmp16 + tmp17;
    assign tans_18_19 = tmp18 + tmp19;
    assign tans_20_21 = tmp20 + tmp21;
    assign tans_22_23 = tmp22 + tmp23;
    assign tans_24_25 = tmp24 + tmp25;
    assign tans_26_27 = tmp26 + tmp27;
    assign tans_28_29 = tmp28 + tmp29;
    assign tans_30_31 = tmp30 + tmp31;
   
    assign tans_01_23 = tans_0_1 + tans_2_3;
    assign tans_45_67 = tans_4_5 + tans_6_7;
    assign tans_89_1011 = tans_8_9 + tans_10_11;
    assign tans_1213_1415 = tans_12_13 + tans_14_15;
    assign tans_1617_1819 = tans_16_17 + tans_18_19;
    assign tans_2021_2223 = tans_20_21 + tans_22_23;
    assign tans_2425_2627 = tans_24_25 + tans_26_27;
    assign tans_2829_3031 = tans_28_29 + tans_30_31;
    
    assign tans_0123_4567 = tans_01_23 + tans_45_67;
    assign tans_891011_12131415 = tans_89_1011 + tans_1213_1415;
    assign tans_16171819_20212223 = tans_1617_1819 + tans_2021_2223;
    assign tans_24252627_28293031 = tans_2425_2627 + tans_2829_3031;
    
    assign tans_012345678_9101112131415 = tans_0123_4567 + tans_891011_12131415;
    assign tans_1617181920212223_2425262728293031 = tans_16171819_20212223 + tans_24252627_28293031;
    
    assign z = tans_012345678_9101112131415 + tans_1617181920212223_2425262728293031;
    
    always @(*)
    begin
        if(reset == 0)
        begin
            tmp0 <= 'b0; tmp1 <= 'b0; tmp2 <= 'b0; tmp3 <= 'b0;
            tmp4 <= 'b0; tmp5 <= 'b0; tmp6 <= 'b0; tmp7 <= 'b0;
            tmp8 <= 'b0; tmp9 <= 'b0; tmp10 <= 'b0; tmp11 <= 'b0;
            tmp12 <= 'b0; tmp13 <= 'b0; tmp14 <= 'b0; tmp15 <= 'b0;
            tmp16 <= 'b0; tmp17 <= 'b0; tmp18 <= 'b0; tmp19 <= 'b0;
            tmp20 <= 'b0; tmp21 <= 'b0; tmp22 <= 'b0; tmp23 <= 'b0;
            tmp24 <= 'b0; tmp25 <= 'b0; tmp26 <= 'b0; tmp27 <= 'b0;
            tmp28 <= 'b0; tmp29 <= 'b0; tmp30 <= 'b0; tmp31 <= 'b0;
        end
        else
        begin
            tmp0 <= b[0] ? {32'b0, a} : 'b0;
            tmp1 <= b[1] ? {31'b0, a, 1'b0} : 'b0;
            tmp2 <= b[2] ? {30'b0, a, 2'b0} : 'b0;
            tmp3 <= b[3] ? {29'b0, a, 3'b0} : 'b0;
            tmp4 <= b[4] ? {28'b0, a, 4'b0} : 'b0;
            tmp5 <= b[5] ? {27'b0, a, 5'b0} : 'b0;
            tmp6 <= b[6] ? {26'b0, a, 6'b0} : 'b0;
            tmp7 <= b[7] ? {25'b0, a, 7'b0} : 'b0;
            tmp8 <= b[8] ? {24'b0, a, 8'b0} : 'b0;
            tmp9 <= b[9] ? {23'b0, a, 9'b0} : 'b0;
            tmp10 <= b[10] ? {22'b0, a, 10'b0} : 'b0;
            tmp11 <= b[11] ? {21'b0, a, 11'b0} : 'b0;
            tmp12 <= b[12] ? {20'b0, a, 12'b0} : 'b0;
            tmp13 <= b[13] ? {19'b0, a, 13'b0} : 'b0;
            tmp14 <= b[14] ? {18'b0, a, 14'b0} : 'b0;
            tmp15 <= b[15] ? {17'b0, a, 15'b0} : 'b0;
            tmp16 <= b[16] ? {16'b0, a, 16'b0} : 'b0;
            tmp17 <= b[17] ? {15'b0, a, 17'b0} : 'b0;
            tmp18 <= b[18] ? {14'b0, a, 18'b0} : 'b0;
            tmp19 <= b[19] ? {13'b0, a, 19'b0} : 'b0;
            tmp20 <= b[20] ? {12'b0, a, 20'b0} : 'b0;
            tmp21 <= b[21] ? {11'b0, a, 21'b0} : 'b0;
            tmp22 <= b[22] ? {10'b0, a, 22'b0} : 'b0;
            tmp23 <= b[23] ? {9'b0, a, 23'b0} : 'b0;
            tmp24 <= b[24] ? {8'b0, a, 24'b0} : 'b0;
            tmp25 <= b[25] ? {7'b0, a, 25'b0} : 'b0;
            tmp26 <= b[26] ? {6'b0, a, 26'b0} : 'b0;
            tmp27 <= b[27] ? {5'b0, a, 27'b0} : 'b0;
            tmp28 <= b[28] ? {4'b0, a, 28'b0} : 'b0;
            tmp29 <= b[29] ? {3'b0, a, 29'b0} : 'b0;
            tmp30 <= b[30] ? {2'b0, a, 30'b0} : 'b0;
            tmp31 <= b[31] ? {1'b0, a, 31'b0} : 'b0;
        end
    end
endmodule
